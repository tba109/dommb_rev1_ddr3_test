
module altclkctrl (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
